module graph

// A node that contains a value of type `T` in the mutable field`val`.
// Nodes are stored on the heap to ensure stable references to them.
@[heap]
pub struct Node[T] {
pub mut:
	val T
}

// An edge contains two references to nodes of type `T` and an integer weight.
@[heap]
pub struct Edge[T] {
pub:
	node1 &Node[T]
	node2 &Node[T]
pub mut:
	weight int = 1
}

pub fn (gr Graph[T]) get_edge[T](node1 &Node[T], node2 &Node[T]) !&Edge[T] {
	if node1 !in gr.adjacency {
		return error('${node1} does not exist')
	}

	return unsafe { gr.adjacency[node1] }[node2] or {
		return error('There exists no edge between ${node1} and ${node2}')
	}
}

// A graph is a list of references to nodes and a list of references to edges made up of these nodes.
// In addition, it holds an adjacency mapping, the keys are the nodes.
// The values are maps where its keys are nodes adjacent to the original node with value
// the index of the edge between these adjacent nodes in the edges list of the graph.
// The field degrees maps the index of a node in the nodes list to the degree of that node.
@[noinit]
pub struct Graph[T] {
	adjacency map[voidptr]map[voidptr]&Edge[T]
pub:
	nodes []&Node[T]
	edges []&Edge[T]
}

// Factory function to create an Graph from a list of nodes
// and a list of edges containing these nodes.
pub fn Graph.create[T](nodes []&Node[T], edges []&Edge[T]) Graph[T] {
	mut adj := map[voidptr]map[voidptr]&Edge[T]{}

	for edge in edges {
		adj[edge.node1][edge.node2] = edge
		adj[edge.node2][edge.node1] = edge
	}

	return Graph[T]{adj, nodes, edges}
}

// Creates a clone of the graph, changes made in a clone will not affect the original graph.
pub fn (gr Graph[T]) clone[T]() Graph[T] {
	mut nodes := []&Node[T]{cap: gr.nodes.len}
	mut edges := []&Edge[T]{cap: gr.edges.len}

	mut adj := map[voidptr]map[voidptr]&Edge[T]{}
	mut node_to_index := map[voidptr]int{}
	for i in 0 .. gr.nodes.len {
		node := &Node[T]{gr.nodes[i].val}
		node_to_index[gr.nodes[i]] = i
		nodes << node
	}

	for edge in gr.edges {
		new_edge := &Edge[T]{nodes[node_to_index[edge.node1]], nodes[node_to_index[edge.node2]], edge.weight}
		edges << new_edge
		adj[edge.node1][edge.node2] = new_edge
		adj[edge.node2][edge.node1] = new_edge
	}

	return Graph[T]{adj, nodes, edges}
}
