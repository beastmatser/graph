module graph

import math

fn test_properties() {
	cycle4 := cycle_graph(4)
	complete6 := complete_graph(6)
	path50 := path_graph(50)
	large := Graph.from_graph6(r'~?Bys????@?O??@?@?@????????????????C??@???O??????????@????_???O??????CA?K?????C_???O????O??@?G???o?_??G?C??@???B?????W?????C?_???D??????O?????????????????O??????O??????O??????G??????C???????G????????????????K???????g????????S???????`?????????????????????????????????????A_???????????A_??????@A???????_???A????@O?????????@?????G??????_???O????@?????_?????G???A??????G???G?????@???G???????@???O?????C????G??????????K????@????????G???_???????_????A??????G?????_?????C???G???????A???????????@_??????_????????????O??????????????G????????????_???????????G?????????????_????????????C?????????????C????????????_?????????????O????????????????????????????????????????????????????????????????????O??????????_??O?????????????C??????????????A@?????????????@??C????????????A?O?????????????O??O???????????G??G????????????A???C????????????C??G????????????@??O????????????G???O???????????????_???????????????A??????????????C??C????????????????_????????????????@???????????????@??O??????????????O??O??????????????_??G?????????????????AA?????????????????G_????????????????AA??????????????????c?????????????????AG?????????????????CO???????????@???????????????????G???????????????????O??????????????????A?????????????????????????????G???????????????????C????????????????????_???????????????????O????????????????????_???????????????????@??????????????????_??O????????????????O??@?????????????????C???_?????????????????O??C?????????????????C???_?????????????????@???_?????????????????G??@?????????????????C???A?????????????????K?????????????????????C?G??????????????????????__????????????????????@_??????????????????????a??????????????????????W?????????????C?????????????????????????????_??????????????????????????????@_???????????????????A??A??????????????????????GG??????????????????????P??????????????????????C?G??????????????????????GO??????????????????????C?_????????????????????@A????????????????????????I???????????????????????@?C???????????????????????GG???????????????????????_?C??????????????????????????K????????????????????????@?A????????????????????????G_????????????????????????P?????????????????????????@C?????????????????????????a?????????@??????????????????????????A??????????????????????????A??????????????????????????@?????????????????????????????????_????????????????????????????C???????????????????????????O??????????????????????????O???????????????????????????O????????????????????????????????????@C???????????????????????????H???????????????????????????D????????????????????????????`???????????????????????????@A???????????????????????????W???????????????????????????O@????????????????????????????_O???????????????????????????_A????????????????????????????_G???????????????????????????G?O??????????????????????????@A??????????????????????????????????????????????????????????????????????????????O?????????????????????????????@??????????????????????????????O??????????????????????????????????????????????????????????????????C???????????????????????????????G??????????????????????????????@???????????????????????????????_??????????????????????????????C???????????????????????????????O?????????????????????????????????????????@O???????????????????????????????_O??????????????????????????????P???????????????????????????????A@???????????????????????????????OG???????????????????????????????__??????????????????????????????CA??????????????????????????????A@???????????????????????????????O?O????????????????????????????????G?C??????????????????????????????_C????????????????????????????????A?@??????????????????????????????A??_???????????????????????????????C?C????????????????????????????????_?_??????????????????????????????C??_???????????????????????????????@??G??????????????????????????????@?@??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????A??@?????????????????????????????????O?G????????????????????????????????@??O????????????????????????????????A??C????????????????????????????????A??A????????????????????????????????@??@??????????????????????????????????W????????????????????????????????????K????????????????????????????????????E????????????????????????????????????`?????????????????????????????????????Q????????????????????????????????????B??????????????????????????????????????OO????????????????????????????????????A_????????????????????????????????????O_????????????????????????????????????GO????????????????????????????????????OA????????????????????????????????????G@???????????????????????????????O??????????????????????????????????????_??????????????????????????????????????C?????????????????????????????????????????????OO?????????????????????????????????????@G?????????????????????????????????????@@??????????????????????????????????????CC??????????????????????????????????????A_??????????????????????????????????????G_???????????????????????????????????G???????????????????????????????????????A???????????????????????????????????????A?????O??????????????????????????????????????OP???????????????????????????????????????_`???????????????????????????????????????C__??????????????????????????????????????G_O??????????????????????????????????????P?G??????????????????????????????????????AG?') or {
		Graph.create[int]([], [])
	}

	// is_bipartite
	assert cycle4.is_bipartite()
	assert path50.is_bipartite()
	assert large.is_bipartite()

	assert !complete6.is_bipartite()

	// is_acyclic
	assert path50.is_acyclic()

	assert !cycle4.is_acyclic()
	assert !large.is_acyclic()
	assert !complete6.is_acyclic()

	// is_connected
	assert cycle4.is_connected()
	assert path50.is_connected()
	assert large.is_connected()
	assert complete6.is_connected()

	// diameter
	assert cycle4.diameter() == 2
	assert path50.diameter() == 49
	assert large.diameter() == 15
	assert complete6.diameter() == 1

	// radius
	assert cycle4.radius() == 2
	assert path50.radius() == 25
	assert large.radius() == 15
	assert complete6.radius() == 1

	// girth
	assert cycle4.girth() == 4
	assert path50.girth() == -1
	assert large.girth() == 6
	assert complete6.girth() == 3

	// num_spanning_trees
	assert cycle4.num_spanning_trees() == 4
	assert path50.num_spanning_trees() == 1
	assert math.log10(large.num_spanning_trees()) - math.log10(2.904638012179e+87) < 1e-12 // small enough
	assert complete6.num_spanning_trees() == 1296

	// num_triangles
	assert cycle4.num_triangles() == 0
	assert path50.num_triangles() == 0
	assert large.num_triangles() == 0
	assert complete6.num_triangles() == 20

	// degeneracy
	assert cycle4.degeneracy() == 2
	assert path50.degeneracy() == 1
	assert large.degeneracy() == 3
	assert complete6.degeneracy() == 5
}
